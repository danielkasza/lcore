/* LC-3 opcodes. */
package opcodes;
/* ADD instructions. */
localparam [15:0] add_rr  = 16'b0001??????000???;
localparam [15:0] add_imm = 16'b0001??????1?????;
/* AND instructions. */
localparam [15:0] and_rr  = 16'b0101??????000???;
localparam [15:0] and_imm = 16'b0101??????1?????;
/* Jump instructions. */
localparam [15:0] br      = 16'b0000????????????;
localparam [15:0] jmp     = 16'b1100000???000000;
localparam [15:0] jsr     = 16'b01001???????????;
localparam [15:0] jsrr    = 16'b0100000???000000;
/* Load instructions. */
localparam [15:0] ld      = 16'b0010????????????;
localparam [15:0] ldr     = 16'b0110????????????;
localparam [15:0] lea     = 16'b1110????????????;
/* XOR instruction.
 * This replaces the LC-3 standard NOT instruction, while maintaining compatiblity.
 * NOT is the same as XOR with 0xFFFF.
 */
localparam [15:0] xor_rr  = 16'b1001??????000???;
localparam [15:0] xor_imm = 16'b1001??????1?????;
/* Interrupt return. */
localparam [15:0] rti     = 16'b1000000000000000;
/* Store instructions. */
localparam [15:0] st      = 16'b0011????????????;
localparam [15:0] str     = 16'b0111????????????;
/* I/O instructions.
 * These use encoding space that was reserved for LDI and STI.
 */
localparam [15:0] in      = 16'b1010????????????;
localparam [15:0] out     = 16'b1011????????????;
/* Bitshift instructions.
 * These were borrowed from the LC-3b ISA.
 */
localparam [15:0] lshf    = 16'b1101??????00????;
localparam [15:0] rshfl   = 16'b1101??????01????;
localparam [15:0] rshfa   = 16'b1101??????11????;
endpackage